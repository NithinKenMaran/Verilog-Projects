`define ADD 3'b001
`define SUB 3'b010
`define AND 3'b011
`define OR 3'b100
`define XOR 3'b101