module control_unit(
    input clk, reset,
    input [3:0] opcode,
    
)