`define ADD 4'b0001
`define SUB 4'b0010
`define AND 4'b0011
`define OR 4'b0100
`define XOR 4'b0101
`define LDR 4'b0110
`define STOP 4'b1111