`define ADD 4'b0000
`define SUB 4'b0001
`define AND 4'b0010
`define OR 4'b0011
`define XOR 4'b0100

`define LDR 4'b0101
`define LPM 4'b0110
`define STM 4'b0111
