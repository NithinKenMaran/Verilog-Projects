module control_unit(
    input clk
);

    // registers //
    reg [1:0] sreg;
    reg [15:0] r [0:7]; // register file


endmodule